module mesh (
    interface node1_PE_in, node1_PE_out,
    node2_PE_in, node2_PE_out,
    node3_PE_in, node3_PE_out,
    node4_PE_in, node4_PE_out,
    node5_PE_in, node5_PE_out,
    node6_PE_in, node6_PE_out,
    node7_PE_in, node7_PE_out,
    node8_PE_in, node8_PE_out,
    node9_PE_in, node9_PE_out,
    node10_PE_in, node10_PE_out,
    node11_PE_in, node11_PE_out,
    node12_PE_in, node12_PE_out,
    node13_PE_in, node13_PE_out,
    node14_PE_in, node14_PE_out,
    node15_PE_in, node15_PE_out
);
    
endmodule