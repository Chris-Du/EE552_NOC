module mesh (
    interface node1_PE_in, node1_PE_out,
    node2_PE_in, node2_PE_out,
    node3_PE_in, node3_PE_out,
    node4_PE_in, node4_PE_out,
    node5_PE_in, node5_PE_out,
    node6_PE_in, node6_PE_out,
    node7_PE_in, node7_PE_out,
    node8_PE_in, node8_PE_out,
    node9_PE_in, node9_PE_out,
    node10_PE_in, node10_PE_out,
    node11_PE_in, node11_PE_out,
    node12_PE_in, node12_PE_out,
    node13_PE_in, node13_PE_out,
    node14_PE_in, node14_PE_out,
    node15_PE_in, node15_PE_out
);
    
    router node1(
        node1_north_in, node1_north_out,
        node1_south_in, node1_south_out, 
        node1_east_in, node1_east_out, 
        node1_west_in, node1_west_out,
        node1_PE_in, node1_PE_out
    );

    router node2(
        node2_north_in, node2_north_out,
        node2_south_in, node2_south_out, 
        node2_east_in, node2_east_out, 
        node2_west_in, node2_west_out,
        node2_PE_in, node2_PE_out
    );

    router node3(
        node3_north_in, node3_north_out,
        node3_south_in, node3_south_out, 
        node3_east_in, node3_east_out, 
        node3_west_in, node3_west_out,
        node3_PE_in, node3_PE_out
    );

    router node4(
        node4_north_in, node4_north_out,
        node4_south_in, node4_south_out, 
        node4_east_in, node4_east_out, 
        node4_west_in, node4_west_out,
        node4_PE_in, node4_PE_out
    );

    router node5(
        node5_north_in, node5_north_out,
        node5_south_in, node5_south_out, 
        node5_east_in, node5_east_out, 
        node5_west_in, node5_west_out,
        node5_PE_in, node5_PE_out
    );

    router node6(
        node6_north_in, node6_north_out,
        node6_south_in, node6_south_out, 
        node6_east_in, node6_east_out, 
        node6_west_in, node6_west_out,
        node6_PE_in, node6_PE_out
    );

    router node7(
        node7_north_in, node7_north_out,
        node7_south_in, node7_south_out, 
        node7_east_in, node7_east_out, 
        node7_west_in, node7_west_out,
        node7_PE_in, node7_PE_out
    );

    router node8(
        node8_north_in, node8_north_out,
        node8_south_in, node8_south_out, 
        node8_east_in, node8_east_out, 
        node8_west_in, node8_west_out,
        node8_PE_in, node8_PE_out
    );
    
    router node9(
        node9_north_in, node9_north_out,
        node9_south_in, node9_south_out, 
        node9_east_in, node9_east_out, 
        node9_west_in, node9_west_out,
        node9_PE_in, node9_PE_out
    );

    router node10(
        node10_north_in, node10_north_out,
        node10_south_in, node10_south_out, 
        node10_east_in, node10_east_out, 
        node10_west_in, node10_west_out,
        node10_PE_in, node10_PE_out
    );

    router node11(
        node11_north_in, node11_north_out,
        node11_south_in, node11_south_out, 
        node11_east_in, node11_east_out, 
        node11_west_in, node11_west_out,
        node11_PE_in, node11_PE_out
    );

    router node12(
        node12_north_in, node12_north_out,
        node12_south_in, node12_south_out, 
        node12_east_in, node12_east_out, 
        node12_west_in, node12_west_out,
        node12_PE_in, node12_PE_out
    );

    router node13(
        node13_north_in, node13_north_out,
        node13_south_in, node13_south_out, 
        node13_east_in, node13_east_out, 
        node13_west_in, node13_west_out,
        node13_PE_in, node13_PE_out
    );

    router node14(
        node14_north_in, node14_north_out,
        node14_south_in, node14_south_out, 
        node14_east_in, node14_east_out, 
        node14_west_in, node14_west_out,
        node14_PE_in, node14_PE_out
    );

    router node15(
        node15_north_in, node15_north_out,
        node15_south_in, node15_south_out, 
        node15_east_in, node15_east_out, 
        node15_west_in, node15_west_out,
        node15_PE_in, node15_PE_out
    );

endmodule